 module BPM_lut(lookup, scaler);
	input [7:0] lookup;
	output [19:0] scaler;
	
	assign scaler =(lookup == 8'd1)   ? 1000000 :
						(lookup == 8'd2)   ? 500000  :
						(lookup == 8'd3)   ? 333333  :
						(lookup == 8'd4)   ? 250000  :
						(lookup == 8'd5)   ? 200000  :
						(lookup == 8'd6)   ? 166667  :
						(lookup == 8'd7)   ? 142857  :
						(lookup == 8'd8)   ? 125000  :
						(lookup == 8'd9)   ? 111111  :
						(lookup == 8'd10)  ? 100000  :
						(lookup == 8'd11)  ? 90909   :
						(lookup == 8'd12)  ? 83333   : 
						(lookup == 8'd13)  ? 76923   :
						(lookup == 8'd14)  ? 71429   : 
						(lookup == 8'd15)  ? 66667   :
						(lookup == 8'd16)  ? 62500   :

						(lookup == 8'd17)  ? 58824 :
						(lookup == 8'd18)  ? 55556 :
						(lookup == 8'd19)  ? 52632 : 
						(lookup == 8'd20)  ? 50000 :
						(lookup == 8'd21)  ? 47619 : 
						(lookup == 8'd22)  ? 45455 :
						(lookup == 8'd23)  ? 43478 :
						(lookup == 8'd24)  ? 41667 :
						(lookup == 8'd25)  ? 40000 :
						(lookup == 8'd26)  ? 38462 :
						(lookup == 8'd27)  ? 37037 :
						(lookup == 8'd28)  ? 35714 :
						(lookup == 8'd29)  ? 34483 :
						(lookup == 8'd30)  ? 33333 : 
						(lookup == 8'd31)  ? 32258 : 
						(lookup == 8'd32)  ? 31250 :

						(lookup == 8'd33)  ? 30303 :
						(lookup == 8'd34)  ? 29412 :
						(lookup == 8'd35)  ? 28571 :
						(lookup == 8'd36)  ? 27778 :
						(lookup == 8'd37)  ? 27027 :
						(lookup == 8'd38)  ? 26316 :
						(lookup == 8'd39)  ? 25641 :
						(lookup == 8'd40)  ? 25000 :
						(lookup == 8'd41)  ? 24390 :
						(lookup == 8'd42)  ? 23810 :
						(lookup == 8'd43)  ? 23256 :
						(lookup == 8'd44)  ? 22727 :
						(lookup == 8'd45)  ? 22222 :
						(lookup == 8'd46)  ? 21739 :
						(lookup == 8'd47)  ? 21277 :
						(lookup == 8'd48)  ? 20833 :

						(lookup == 8'd49)  ? 20408 :
						(lookup == 8'd50)  ? 20000 :
						(lookup == 8'd51)  ? 19608 :
						(lookup == 8'd52)  ? 19231 : 
						(lookup == 8'd53)  ? 18868 :
						(lookup == 8'd54)  ? 18519 : 
						(lookup == 8'd55)  ? 18182 :
						(lookup == 8'd56)  ? 17857 :
						(lookup == 8'd57)  ? 17544 : 
						(lookup == 8'd58)  ? 17241 :
						(lookup == 8'd59)  ? 16949 :
						(lookup == 8'd60)  ? 16667 :
						(lookup == 8'd61)  ? 16393 :
						(lookup == 8'd62)  ? 16129 :
						(lookup == 8'd63)  ? 15873 :
						(lookup == 8'd64)  ? 15625 :

						(lookup == 8'd65)  ? 15385 :
						(lookup == 8'd66)  ? 15152 :
						(lookup == 8'd67)  ? 14925 :
						(lookup == 8'd68)  ? 14706 :
						(lookup == 8'd69)  ? 14493 :
						(lookup == 8'd70)  ? 14286 :
						(lookup == 8'd71)  ? 14085 :
						(lookup == 8'd72)  ? 13889 :
						(lookup == 8'd73)  ? 13699 :
						(lookup == 8'd74)  ? 13514 :
						(lookup == 8'd75)  ? 13333 :
						(lookup == 8'd76)  ? 13158 :
						(lookup == 8'd77)  ? 12987 :
						(lookup == 8'd78)  ? 12821 :
						(lookup == 8'd79)  ? 12658 :
						(lookup == 8'd80)  ? 12500 :

						(lookup == 8'd81)  ? 12346 :
						(lookup == 8'd82)  ? 12195 :
						(lookup == 8'd83)  ? 12048 :
						(lookup == 8'd84)  ? 11905 :
						(lookup == 8'd85)  ? 11765 :
						(lookup == 8'd86)  ? 11628 :
						(lookup == 8'd87)  ? 11494 :
						(lookup == 8'd88)  ? 11364 :
						(lookup == 8'd89)  ? 11236 :
						(lookup == 8'd90)  ? 11111 :
						(lookup == 8'd91)  ? 10989 :
						(lookup == 8'd92)  ? 10870 :
						(lookup == 8'd93)  ? 10753 :
						(lookup == 8'd94)  ? 10638 :
						(lookup == 8'd95)  ? 10526 :
						(lookup == 8'd96)  ? 10417 : 

						(lookup == 8'd97)  ? 10309 :
						(lookup == 8'd98)  ? 10204 :
						(lookup == 8'd99)  ? 10101 :
						(lookup == 8'd100) ? 10000 :
						(lookup == 8'd101) ? 9901 : 
						(lookup == 8'd102) ? 9804 :
						(lookup == 8'd103) ? 9709 :
						(lookup == 8'd104) ? 9615 :
						(lookup == 8'd105) ? 9524 :
						(lookup == 8'd106) ? 9434 :
						(lookup == 8'd107) ? 9346 :
						(lookup == 8'd108) ? 9259 :
						(lookup == 8'd109) ? 9174 :
						(lookup == 8'd110) ? 9091 :
						(lookup == 8'd111) ? 9009 :
						(lookup == 8'd112) ? 8929 :

						(lookup == 8'd113) ? 8850 :
						(lookup == 8'd114) ? 8772 :
						(lookup == 8'd115) ? 8696 :
						(lookup == 8'd116) ? 8621 :
						(lookup == 8'd117) ? 8547 :
						(lookup == 8'd118) ? 8475 :
						(lookup == 8'd119) ? 8403 :
						(lookup == 8'd120) ? 8333 :
						(lookup == 8'd121) ? 8264 :
						(lookup == 8'd122) ? 8197 :
						(lookup == 8'd123) ? 8130 :
						(lookup == 8'd124) ? 8065 :
						(lookup == 8'd125) ? 8000 :
						(lookup == 8'd126) ? 7937 :
						(lookup == 8'd127) ? 7874 :
						(lookup == 8'd128) ? 7813 :

						(lookup == 8'd129) ? 7752 :
						(lookup == 8'd130) ? 7692 :
						(lookup == 8'd131) ? 7634 :
						(lookup == 8'd132) ? 7576 :
						(lookup == 8'd133) ? 7519 :
						(lookup == 8'd134) ? 7463 :
						(lookup == 8'd135) ? 7407 :
						(lookup == 8'd136) ? 7353 :
						(lookup == 8'd137) ? 7299 :
						(lookup == 8'd138) ? 7246 :
						(lookup == 8'd139) ? 7194 : 
						(lookup == 8'd140) ? 7143 :
						(lookup == 8'd141) ? 7092 :
						(lookup == 8'd142) ? 7042 :
						(lookup == 8'd143) ? 6993 :
						(lookup == 8'd144) ? 6944 :

						(lookup == 8'd145) ? 6897 :
						(lookup == 8'd146) ? 6849 :
						(lookup == 8'd147) ? 6803 :
						(lookup == 8'd148) ? 6757 :
						(lookup == 8'd149) ? 6711 :
						(lookup == 8'd150) ? 6667 :
						(lookup == 8'd151) ? 6623 :
						(lookup == 8'd152) ? 6579 :
						(lookup == 8'd153) ? 6536 :
						(lookup == 8'd154) ? 6494 :
						(lookup == 8'd155) ? 6452 :
						(lookup == 8'd156) ? 6410 :
						(lookup == 8'd157) ? 6369 :
						(lookup == 8'd158) ? 6329 :
						(lookup == 8'd159) ? 6289 :
						(lookup == 8'd160) ? 6250 :

						(lookup == 8'd161) ? 6211 :
						(lookup == 8'd162) ? 6173 :
						(lookup == 8'd163) ? 6135 :
						(lookup == 8'd164) ? 6098 :
						(lookup == 8'd165) ? 6061 : 
						(lookup == 8'd166) ? 6024 :
						(lookup == 8'd167) ? 5988 :
						(lookup == 8'd168) ? 5952 :
						(lookup == 8'd169) ? 5917 :
						(lookup == 8'd170) ? 5882 :
						(lookup == 8'd171) ? 5848 :
						(lookup == 8'd172) ? 5814 :
						(lookup == 8'd173) ? 5780 :
						(lookup == 8'd174) ? 5747 :
						(lookup == 8'd175) ? 5714 :
						(lookup == 8'd176) ? 5682 :

						(lookup == 8'd177) ? 5650 :
						(lookup == 8'd178) ? 5618 :
						(lookup == 8'd179) ? 5587 :
						(lookup == 8'd180) ? 5556 :
						(lookup == 8'd181) ? 5525 :
						(lookup == 8'd182) ? 5495 :
						(lookup == 8'd183) ? 5464 :
						(lookup == 8'd184) ? 5435 :
						(lookup == 8'd185) ? 5405 :
						(lookup == 8'd186) ? 5376 :
						(lookup == 8'd187) ? 5348 :
						(lookup == 8'd188) ? 5319 :
						(lookup == 8'd189) ? 5291 :
						(lookup == 8'd190) ? 5263 :
						(lookup == 8'd191) ? 5236 :
						(lookup == 8'd192) ? 5208 :

						(lookup == 8'd193) ? 5181 :
						(lookup == 8'd194) ? 5155 :
						(lookup == 8'd195) ? 5128 : 
						(lookup == 8'd196) ? 5102 :
						(lookup == 8'd197) ? 5076 :
						(lookup == 8'd198) ? 5051 :
						(lookup == 8'd199) ? 5025 :
						(lookup == 8'd200) ? 5000 :
						(lookup == 8'd201) ? 4975 :
						(lookup == 8'd202) ? 4950 :
						(lookup == 8'd203) ? 4926 :
						(lookup == 8'd204) ? 4902 :
						(lookup == 8'd205) ? 4878 :
						(lookup == 8'd206) ? 4854 :
						(lookup == 8'd207) ? 4831 :
						(lookup == 8'd208) ? 4808 :

						(lookup == 8'd209) ? 4785 :
						(lookup == 8'd210) ? 4762 :
						(lookup == 8'd211) ? 4739 :
						(lookup == 8'd212) ? 4717 :
						(lookup == 8'd213) ? 4695 :
						(lookup == 8'd214) ? 4673 :
						(lookup == 8'd215) ? 4651 :
						(lookup == 8'd216) ? 4630 :
						(lookup == 8'd217) ? 4608 :
						(lookup == 8'd218) ? 4587 :
						(lookup == 8'd219) ? 4566 :
						(lookup == 8'd220) ? 4545 :
						(lookup == 8'd221) ? 4525 : 
						(lookup == 8'd222) ? 4505 :
						(lookup == 8'd223) ? 4484 :
						(lookup == 8'd224) ? 4464 :

						(lookup == 8'd225) ? 4444 :
						(lookup == 8'd226) ? 4425 :
						(lookup == 8'd227) ? 4405 :
						(lookup == 8'd228) ? 4386 :
						(lookup == 8'd229) ? 4367 :
						(lookup == 8'd230) ? 4348 :
						(lookup == 8'd231) ? 4329 :
						(lookup == 8'd232) ? 4310 :
						(lookup == 8'd233) ? 4292 :
						(lookup == 8'd234) ? 4274 :
						(lookup == 8'd235) ? 4255 :
						(lookup == 8'd236) ? 4237 :
						(lookup == 8'd237) ? 4219 :
						(lookup == 8'd238) ? 4202 :
						(lookup == 8'd239) ? 4184 :
						(lookup == 8'd240) ? 4167 :

						(lookup == 8'd241) ? 4149 :
						(lookup == 8'd242) ? 4132 :
						(lookup == 8'd243) ? 4115 :
						(lookup == 8'd244) ? 4098 :
						(lookup == 8'd245) ? 4082 :
						(lookup == 8'd246) ? 4065 :
						(lookup == 8'd247) ? 4049 :
						(lookup == 8'd248) ? 4032 : 
						(lookup == 8'd249) ? 4016 :
						(lookup == 8'd250) ? 4000 :
						(lookup == 8'd251) ? 3984 :
						(lookup == 8'd252) ? 3968 :
						(lookup == 8'd253) ? 3953 :
						(lookup == 8'd254) ? 3937 :
						(lookup == 8'd255) ? 3922 :
						/*lookup undef*/ 20'hFFFFF;

endmodule
